`timescale 1ns / 1ps



module tb_Asynchronous_RAM_port1(

    );
endmodule
